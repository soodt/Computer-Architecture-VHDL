library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- Uncomment the following library declaration if using-- arithmetic functions with Signed or Unsigned architectureuse IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if instantiating-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
entity CPU_ControlMemory_21356526 is
	Port ( Address : in STD_LOGIC_VECTOR (16 downto 0);
		  NA : out STD_LOGIC_VECTOR (16 downto 0); -- 34-50
		  MS : out STD_LOGIC_VECTOR (2 downto 0); -- 31-33
		MC : out STD_LOGIC; -- 30
		IL : out STD_LOGIC; -- 29
		PI : out STD_LOGIC; -- 28
		PL : out STD_LOGIC; -- 27
		TD : out STD_LOGIC_VECTOR (3 downto 0); -- 23-26
		TA : out STD_LOGIC_VECTOR (3 downto 0); -- 19-22
		TB : out STD_LOGIC_VECTOR (3 downto 0); -- 15-18
		MB : out STD_LOGIC; -- 14
		FS : out STD_LOGIC_VECTOR (4 downto 0); -- 09-13
		MD : out STD_LOGIC; -- 08
		RW : out STD_LOGIC; -- 07
		MM : out STD_LOGIC; -- 06
		MW : out STD_LOGIC; -- 05
		RV : out STD_LOGIC; -- 04
		RC : out STD_LOGIC; -- 03
		RN : out STD_LOGIC; -- 02
		RZ : out STD_LOGIC; -- 01
		FL : out STD_LOGIC); -- 00 
end CPU_ControlMemory_21356526;
architecture Behavioral of CPU_ControlMemory_21356526 is
-- we use the least significant 7 bit of the Address - array(0 to 127)
type ROM_array is array(0 to 127) of STD_LOGIC_VECTOR (50 downto 0);
signal ROM : ROM_array :=(
--|50               34|33 31| 30| 29| 28| 27|26 23|22 19  |18 15 | 14|13   09| 08| 07| 06| 05| 04| 03| 02| 01| 00| Control Mem     s
--| Next Address      |  MS | MC| IL| PI| PL| TD  | TA    |  TB  | MB| FS    | MD| RW| MM| MW| RV| RC| RN| RZ| FL| Address
   "00000000000000000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 00
   "00000000000000001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 01
   "00000000000000010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 02
   "00000000000000011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 03
   "00000000000000100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 04
   "00000000000000101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 05       
   "00000000000000110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 06  
   "00000000000000111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 07  
   "00000000000001000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 08
   "00000000000001001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 09  
   "00000000000001010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 0A  
   "00000000000001011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 0B  
   "00000000000001100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 0C 
   "00000000000001101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 0D 
   "00000000000001110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 0E 
   "00000000000001111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 0F
   "00000000000010001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 11     "00000000000010010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 12 "00000000000010011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 13 "00000000000010100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 14 "00000000000010101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 15 "00000000000010110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 16 "00000000000010111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 17 "00000000000011000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 18 "00000000000011001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 19 "00000000000011010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 1A "00000000000011011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 1B "00000000000011100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 1C "00000000000011101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 1D "00000000000011110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 1E "00000000000011111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 1F 
   "00000000001110000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 70
   "00000000001110001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 71
   "00000000001110010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 72
   "00000000001110011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 73
   "00000000001110100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 74
   "00000000001110101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 75
   "00000000001110110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 76
   "00000000001110111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 77
   "00000000001111000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 78
   "00000000001111001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 79
   "00000000001111010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 7A
   "00000000001111011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 7B
   "00000000001111100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 7C
   "00000000001111101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 7D
   "00000000001111110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0', -- 7E
   "00000000001111111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0' -- 7F 
);

signal content_at_address : STD_LOGIC_VECTOR (50 downto 0); 

begin
content_at_address <= ROM(to_integer(unsigned(Address(6 downto 0)))) after 2ns;
NA <= content_at_address(50 downto 34); -- 34-50
MS <= content_at_address(33 downto 31);  -- 31-33
MC <= content_at_address(30);            -- 30
IL <= content_at_address(29);            -- 29
PI <= content_at_address(28);            -- 28
PL <= content_at_address(27);            -- 27
TD <= content_at_address(26 downto 23);  -- 23-26
TA <= content_at_address(22 downto 19);  -- 19-22
TB <= content_at_address(18 downto 15);  -- 15-18
MB <= content_at_address(14); 		 -- 14
FS <= content_at_address(13 downto 9);   -- 09-13
MD <= content_at_address(8); 		 -- 08
RW <= content_at_address(7); 		 -- 07
MM <= content_at_address(6); 		 -- 06
MW <= content_at_address(5); 		 -- 05
RV <= content_at_address(4); 		 -- 04
RC <= content_at_address(3); 		 -- 03
RN <= content_at_address(2); 		 -- 02
RZ <= content_at_address(1); 		 -- 01
FL <= content_at_address(0);		 -- 00
end Behavioral;
