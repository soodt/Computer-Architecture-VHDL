library ieee; 
use ieee.std_logic_1164.all; 
entity DP_RippleCarryAdder32Bit_21356526 is
port(B, A : in std_logic_vector(31 downto 0);
 	C_IN: in std_logic; 
	SUM : out std_logic_vector(31 downto 0); 
	C_OUT : out std_logic; 
	V : out STD_LOGIC);
end DP_RippleCarryAdder32Bit_21356526;

architecture Behavioral of DP_RippleCarryAdder32Bit_21356526 is

COMPONENT DP_FullAdder_21356526   
    PORT(
         A : in STD_LOGIC;
         B : in STD_LOGIC;
         C_IN : in STD_LOGIC;
         SUM : out STD_LOGIC;
         C_OUT : out STD_LOGIC
        );
END COMPONENT;

Signal C0,  C1,  C2,  C3,  C4,  C5,  C6,  C7,  C8,  C9,  C10,  C11,  C12,  C13,  C14,  C15,  C16,  C17,  C18,  C19,  C20,  C21,  C22,  C23,  C24,  C25,  C26,  C27,  C28,  C29,  C30,  C31 : STD_LOGIC;

begin

BIT0: DP_FullAdder_21356526 PORT MAP (
       A => A(0),
       B => B(0),
       C_IN => C_IN,
       SUM => SUM(0),
       C_OUT => C0
      );
BIT1: DP_FullAdder_21356526 PORT MAP (
       A => A(1),
       B => B(1),
       C_IN => C0,
       SUM => SUM(1),
       C_OUT => C1
      );
BIT2: DP_FullAdder_21356526 PORT MAP (
       A => A(2),
       B => B(2),
       C_IN => C1,
       SUM => SUM(2),
       C_OUT => C2
      );
BIT3: DP_FullAdder_21356526 PORT MAP (
       A => A(3),
       B => B(3),
       C_IN => C2,
       SUM => SUM(3),
       C_OUT => C3
      );
BIT4: DP_FullAdder_21356526 PORT MAP (
       A => A(4),
       B => B(4),
       C_IN => C3,
       SUM => SUM(4),
       C_OUT => C4
      );
BIT5: DP_FullAdder_21356526 PORT MAP (
       A => A(5),
       B => B(5),
       C_IN => C4,
       SUM => SUM(5),
       C_OUT => C5
      );
BIT6: DP_FullAdder_21356526 PORT MAP (
       A => A(6),
       B => B(6),
       C_IN => C5,
       SUM => SUM(6),
       C_OUT => C6
      );
BIT7: DP_FullAdder_21356526 PORT MAP (
       A => A(7),
       B => B(7),
       C_IN => C6,
       SUM => SUM(7),
       C_OUT => C7
      );
BIT8: DP_FullAdder_21356526 PORT MAP (
       A => A(8),
       B => B(8),
       C_IN => C7,
       SUM => SUM(8),
       C_OUT => C8
      );
BIT9: DP_FullAdder_21356526 PORT MAP (
       A => A(9),
       B => B(9),
       C_IN => C8,
       SUM => SUM(9),
       C_OUT => C9
      );
BIT10: DP_FullAdder_21356526 PORT MAP (
       A => A(10),
       B => B(10),
       C_IN => C9,
       SUM => SUM(10),
       C_OUT => C10
      );
BIT11: DP_FullAdder_21356526 PORT MAP (
       A => A(11),
       B => B(11),
       C_IN => C10,
       SUM => SUM(11),
       C_OUT => C11
      );
BIT12: DP_FullAdder_21356526 PORT MAP (
       A => A(12),
       B => B(12),
       C_IN => C11,
       SUM => SUM(12),
       C_OUT => C12
      );
BIT13: DP_FullAdder_21356526 PORT MAP (
       A => A(13),
       B => B(13),
       C_IN => C12,
       SUM => SUM(13),
       C_OUT => C13
      );
BIT14: DP_FullAdder_21356526 PORT MAP (
       A => A(14),
       B => B(14),
       C_IN => C13,
       SUM => SUM(14),
       C_OUT => C14
      );
BIT15: DP_FullAdder_21356526 PORT MAP (
       A => A(15),
       B => B(15),
       C_IN => C14,
       SUM => SUM(15),
       C_OUT => C15
      );
BIT16: DP_FullAdder_21356526 PORT MAP (
       A => A(16),
       B => B(16),
       C_IN => C15,
       SUM => SUM(16),
       C_OUT => C16
      );
BIT17: DP_FullAdder_21356526 PORT MAP (
       A => A(17),
       B => B(17),
       C_IN => C16,
       SUM => SUM(17),
       C_OUT => C17
      );
BIT18: DP_FullAdder_21356526 PORT MAP (
       A => A(18),
       B => B(18),
       C_IN => C17,
       SUM => SUM(18),
       C_OUT => C18
      );
BIT19: DP_FullAdder_21356526 PORT MAP (
       A => A(19),
       B => B(19),
       C_IN => C18,
       SUM => SUM(19),
       C_OUT => C19
      );
BIT20: DP_FullAdder_21356526 PORT MAP (
       A => A(20),
       B => B(20),
       C_IN => C19,
       SUM => SUM(20),
       C_OUT => C20
      );
BIT21: DP_FullAdder_21356526 PORT MAP (
       A => A(21),
       B => B(21),
       C_IN => C20,
       SUM => SUM(21),
       C_OUT => C21
      );
BIT22: DP_FullAdder_21356526 PORT MAP (
       A => A(22),
       B => B(22),
       C_IN => C21,
       SUM => SUM(22),
       C_OUT => C22
      );
BIT23: DP_FullAdder_21356526 PORT MAP (
       A => A(23),
       B => B(23),
       C_IN => C22,
       SUM => SUM(23),
       C_OUT => C23
      );
BIT24: DP_FullAdder_21356526 PORT MAP (
       A => A(24),
       B => B(24),
       C_IN => C23,
       SUM => SUM(24),
       C_OUT => C24
      );
BIT25: DP_FullAdder_21356526 PORT MAP (
       A => A(25),
       B => B(25),
       C_IN => C24,
       SUM => SUM(25),
       C_OUT => C25
      );
BIT26: DP_FullAdder_21356526 PORT MAP (
       A => A(26),
       B => B(26),
       C_IN => C25,
       SUM => SUM(26),
       C_OUT => C26
      );
BIT27: DP_FullAdder_21356526 PORT MAP (
       A => A(27),
       B => B(27),
       C_IN => C26,
       SUM => SUM(27),
       C_OUT => C27
      );
BIT28: DP_FullAdder_21356526 PORT MAP (
       A => A(28),
       B => B(28),
       C_IN => C27,
       SUM => SUM(28),
       C_OUT => C28
      );
BIT29: DP_FullAdder_21356526 PORT MAP (
       A => A(29),
       B => B(29),
       C_IN => C28,
       SUM => SUM(29),
       C_OUT => C29
      );
BIT30: DP_FullAdder_21356526 PORT MAP (
       A => A(30),
       B => B(30),
       C_IN => C29,
       SUM => SUM(30),
       C_OUT => C30
      );
BIT31: DP_FullAdder_21356526 PORT MAP (
       A => A(31),
       B => B(31),
       C_IN => C30,
       SUM => SUM(31),
       C_OUT => C31
      );

C_OUT <= C31;
V <= C31 XOR C1 after 3ns;

end Behavioral;
